module top(
    input               clk,
    input               rst_n,

    output reg [3:0]    led = 4'b0001
);

parameter CLK_FRE = 50;

/********************************************************************************/
/**************************    计数器分频    ************************************/
/********************************************************************************/
reg [31:0] cnt = 0;
always@(posedge clk or negedge rst_n) 
    if(!rst_n) 
        cnt <= 0;
    else 
        cnt <= (cnt >= CLK_FRE * 1000_000 -1)? 0: cnt + 1;

/********************************************************************************/
/**************************     移位显示    ************************************/
/********************************************************************************/
always@(posedge clk or negedge rst_n) 
    if(!rst_n) 
        led <= 4'b0001;
    else 
        if(cnt == 0)
            led <= {led[2:0], led[3]};
        else 
            led <= led;

endmodule